`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:01:00 04/23/2015 
// Design Name: 
// Module Name:    modBigNumbers 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module modBigNumbers(
    input [63:0] exponent,
    input [63:0] number,
    input [63:0] logNum,
    output reg [31:0] result
    );
	 
	 


endmodule
